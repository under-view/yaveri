ADed_$;
_fea9213;
shiftreg_a;
busa_index;
error_condition;
merge_ab;
_bus3;
n$657;
