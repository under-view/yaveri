ADed_$;
_fea9213;
9dae;
$dae;
