\busa+index
\-clock
\***error-condition***
\net1/\net2
\{a,b}
\a*(b+c)
\net           // "net" is a keyword. "\net " is a user-defined identifier.
