\busa+index
\-clock
\***error-condition***
\net1/\net2
\{a,b}
\a*(b+c)
\net
