// this file should not generate any output
// here is a comment
/* here is a simple comment */
/* here 
is 
a 
multi-line
comment
*/

/* here are some nasty comments: */
/* ///// /// */
/*******/
