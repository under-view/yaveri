$display ("display a message");
$finish;
